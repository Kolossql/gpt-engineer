module lfsr_tb;

  reg clk;
  reg reset;
  wire [7:0] data;

  lfsr uut (
    .clk(clk),
    .reset(reset),
    .data(data)
  );

  always begin
    #5 clk = ~clk;
  end

  initial begin
    clk = 0;
    reset = 1;
    #10 reset = 0;
    #100 $finish;
  end

endmodule
